*** SPICE deck for cell xor-gate{lay} from library xor-gate
*** Created on Mon Sep 25, 2023 20:41:36
*** Last revised on Wed Sep 27, 2023 19:29:06
*** Written on Wed Sep 27, 2023 19:34:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: xor-gate{lay}
Mnmos@0 net@1 A gnd gnd N L=0.35U W=1.4U AS=4.563P AD=1.593P PS=11.681U PD=5.075U
Mnmos@1 net@3 B gnd gnd N L=0.35U W=1.4U AS=4.563P AD=1.593P PS=11.681U PD=5.075U
Mnmos@2 F B net@14 gnd N L=0.35U W=1.4U AS=1.378P AD=1.348P PS=4.069U PD=4.025U
Mnmos@3 net@14 net@1 F gnd N L=0.35U W=1.4U AS=1.348P AD=1.378P PS=4.025U PD=4.069U
Mnmos@4 gnd A net@14 gnd N L=0.35U W=1.4U AS=1.378P AD=4.563P PS=4.069U PD=11.681U
Mnmos@5 net@14 net@3 gnd gnd N L=0.35U W=1.4U AS=4.563P AD=1.378P PS=11.681U PD=4.069U
Mpmos@0 net@5 B F vdd P L=0.35U W=1.4U AS=1.348P AD=0.513P PS=4.025U PD=2.188U
Mpmos@1 vdd net@1 net@5 vdd P L=0.35U W=1.4U AS=0.513P AD=4.563P PS=2.188U PD=10.675U
Mpmos@2 net@8 A vdd vdd P L=0.35U W=1.4U AS=4.563P AD=0.482P PS=10.675U PD=2.363U
Mpmos@3 F net@3 net@8 vdd P L=0.35U W=1.4U AS=0.482P AD=1.348P PS=2.363U PD=4.025U
Mpmos@4 net@3 B vdd vdd P L=0.35U W=1.4U AS=4.563P AD=1.593P PS=10.675U PD=5.075U
Mpmos@5 net@1 A vdd vdd P L=0.35U W=1.4U AS=4.563P AD=1.593P PS=10.675U PD=5.075U

* Spice Code nodes in cell cell 'xor-gate{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
VA A 0 PULSE(3.3 0 0 2n 3n 250n 500n)
VB B 0 PULSE(3.3 0 0 2n 3n 125n 250n)
.TRAN 0 1000n
.include Z:\MOS_model.txt
.END
