*** SPICE deck for cell 2to1-mux-schematic{sch} from library 2to1-mux
*** Created on Wed Oct 25, 2023 17:18:56
*** Last revised on Wed Oct 25, 2023 18:14:56
*** Written on Wed Oct 25, 2023 18:15:01 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 2to1-mux-schematic{sch}
Mnmos@0 net@40 S gnd gnd N L=0.35U W=1.4U
Mnmos@1 net@11 net@40 gnd gnd N L=0.35U W=1.4U
Mnmos@2 net@12 S gnd gnd N L=0.35U W=1.4U
Mnmos@3 net@13 D0 net@11 gnd N L=0.35U W=1.4U
Mnmos@4 net@13 D1 net@12 gnd N L=0.35U W=1.4U
Mnmos@5 Y net@13 gnd gnd N L=0.35U W=1.4U
Mpmos@0 net@40 S vdd vdd P L=0.35U W=1.4U
Mpmos@1 net@13 S net@24 vdd P L=0.35U W=1.4U
Mpmos@2 net@13 D1 net@24 vdd P L=0.35U W=1.4U
Mpmos@3 net@24 net@40 vdd vdd P L=0.35U W=1.4U
Mpmos@4 net@24 D0 vdd vdd P L=0.35U W=1.4U
Mpmos@5 Y net@13 vdd vdd P L=0.35U W=1.4U

* Spice Code nodes in cell cell '2to1-mux-schematic{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
*
VS S 0 PULSE(3.3 0 0 1n 1n 500n 1000n)
VD0 D0 0 PULSE(3.3 0 0 1n 1n 100n 200n)
VD1 D1 0 PULSE(3.3 0 0 1n 1n 50n 100n)
*
.TRAN 0 2000n
.include Z:\MOS_model.txt
.END
