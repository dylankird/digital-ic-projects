*** SPICE deck for cell xor-gate{sch} from library xor-gate
*** Created on Mon Sep 25, 2023 17:08:15
*** Last revised on Fri Sep 29, 2023 13:28:28
*** Written on Fri Sep 29, 2023 13:40:04 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: xor-gate{sch}
Mnmos@0 net@83 B gnd gnd N L=0.35U W=1.4U
Mnmos@1 net@62 A gnd gnd N L=0.35U W=1.4U
Mnmos@2 F net@62 net@64 gnd N L=0.35U W=1.4U
Mnmos@3 F B net@64 gnd N L=0.35U W=1.4U
Mnmos@4 net@64 A gnd gnd N L=0.35U W=1.4U
Mnmos@5 net@64 net@83 gnd gnd N L=0.35U W=1.4U
Mpmos@0 net@83 B vdd vdd P L=0.35U W=1.4U
Mpmos@1 net@62 A vdd vdd P L=0.35U W=1.4U
Mpmos@2 net@31 net@62 vdd vdd P L=0.35U W=1.4U
Mpmos@3 F B net@31 vdd P L=0.35U W=1.4U
Mpmos@4 net@19 A vdd vdd P L=0.35U W=1.4U
Mpmos@5 F net@83 net@19 vdd P L=0.35U W=1.4U

* Spice Code nodes in cell cell 'xor-gate{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
*
*For logic simulation:
VA A 0 PULSE(3.3 0 0 2n 3n 250n 500n)
VB B 0 PULSE(3.3 0 0 2n 3n 125n 250n)
*
*For measurements:
*VA A 0 DC 3.3
*VB B 0 PULSE(3.3 0 0 100p 100p 125n 250n)
*
.TRAN 0 1000n
.meas risetime TRIG v(F)=0.33 TD=0 rise=1 TARG v(F)=2.97 TD=0 rise=1
.meas falltime TRIG v(F)=2.97 TD=0 fall=1 TARG v(F)=0.33 TD=0 fall=1
.meas tpHL TRIG v(B)=1.65 TD=0 rise=1 TARG v(F)=1.65 TD=0 fall=1
.meas tpLH TRIG v(B)=1.65 TD=0 fall=1 TARG v(F)=1.65 TD=0 rise=1
.meas propagationdelay param=(tpHL+tpLH)/2
.include Z:\MOS_model.txt
.END
