*** SPICE deck for cell hw3-function-layout{lay} from library hw3-function
*** Created on Mon Nov 06, 2023 10:55:00
*** Last revised on Mon Nov 06, 2023 22:20:06
*** Written on Mon Nov 06, 2023 22:20:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: hw3-function-layout{lay}
Mnmos@1 F X net@7 gnd N L=0.35U W=1.4U AS=0.98P AD=1.593P PS=2.8U PD=5.075U
Mnmos@2 net@7 Z net@9 gnd N L=0.35U W=1.4U AS=0.98P AD=0.98P PS=2.8U PD=2.8U
Mnmos@4 net@7 W net@9 gnd N L=0.35U W=1.4U AS=0.98P AD=0.98P PS=2.8U PD=2.8U
Mnmos@5 net@9 CLK gnd gnd N L=0.35U W=1.4U AS=13.077P AD=0.98P PS=33.075U PD=2.8U
Mnmos@6 net@9 Y net@7 gnd N L=0.35U W=1.4U AS=0.98P AD=0.98P PS=2.8U PD=2.8U
Mpmos@0 F CLK vdd vdd P L=0.35U W=1.4U AS=15.374P AD=1.593P PS=33.425U PD=5.075U

* Spice Code nodes in cell cell 'hw3-function-layout{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
*
*For logic simulation:
VW W 0 PULSE(3.3 0 0 1n 1n 1000n 2000n)
VX X 0 PULSE(3.3 0 0 1n 1n 500n 1000n)
VY Y 0 PULSE(3.3 0 0 1n 1n 250n 500n)
VZ Z 0 PULSE(3.3 0 0 1n 1n 125n 250n)
VCLK CLK 0 PULSE(3.3 0 0 1n 1n 62.5n 125n)
*
.TRAN 0 2000n
.include Z:\MOS_model.txt
.END
