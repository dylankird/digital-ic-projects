*** SPICE deck for cell 8to1-mux-cmos-layout{lay} from library 8to1-mux-cmos
*** Created on Thu Oct 26, 2023 18:37:36
*** Last revised on Thu Oct 26, 2023 20:02:11
*** Written on Thu Oct 26, 2023 20:02:16 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: 8to1-mux-cmos:8to1-mux-cmos-layout{lay}
Mnmos@5 gnd net@141 net@112 gnd N L=0.35U W=1.4U AS=1.593P AD=1.184P PS=5.075U PD=3.558U
Mnmos@6 net@132 S gnd gnd N L=0.35U W=1.4U AS=1.184P AD=0.482P PS=3.558U PD=2.363U
Mnmos@7 Y D1 net@132 gnd N L=0.35U W=1.4U AS=0.482P AD=0.98P PS=2.363U PD=2.8U
Mnmos@8 net@112 D0 Y gnd N L=0.35U W=1.4U AS=0.98P AD=1.593P PS=2.8U PD=5.075U
Mnmos@9 net@141 S gnd gnd N L=0.35U W=1.4U AS=1.184P AD=1.593P PS=3.558U PD=5.075U
Mpmos@5 net@105 net@141 vdd vdd P L=0.35U W=1.4U AS=1.593P AD=0.98P PS=5.075U PD=2.8U
Mpmos@6 Y S net@105 vdd P L=0.35U W=1.4U AS=0.98P AD=0.98P PS=2.8U PD=2.8U
Mpmos@7 net@105 D1 Y vdd P L=0.35U W=1.4U AS=0.98P AD=0.98P PS=2.8U PD=2.8U
Mpmos@8 vdd D0 net@105 vdd P L=0.35U W=1.4U AS=0.98P AD=1.593P PS=2.8U PD=5.075U
Mpmos@9 net@141 S vdd vdd P L=0.35U W=1.4U AS=1.593P AD=1.593P PS=5.075U PD=5.075U

* Spice Code nodes in cell cell '8to1-mux-cmos:8to1-mux-cmos-layout{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
*
VS S 0 PULSE(3.3 0 0 1n 1n 500n 1000n)
VD0 D0 0 PULSE(3.3 0 0 1n 1n 100n 200n)
VD1 D1 0 PULSE(3.3 0 0 1n 1n 50n 100n)
*
.TRAN 0 2000n
.include Z:\MOS_model.txt
.END
