*** SPICE deck for cell 2-input-nand-schematic{sch} from library 2-input-nand
*** Created on Wed Nov 29, 2023 13:23:46
*** Last revised on Wed Nov 29, 2023 18:16:59
*** Written on Wed Nov 29, 2023 18:17:59 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 2-input-nand:2-input-nand-schematic{sch}
Mnmos@0 F A net@0 gnd N L=0.35U W=1.4U
Mnmos@1 net@0 B gnd gnd N L=0.35U W=1.4U
Mpmos@0 F A vdd vdd P L=0.35U W=1.4U
Mpmos@1 F B vdd vdd P L=0.35U W=1.4U

* Spice Code nodes in cell cell '2-input-nand:2-input-nand-schematic{sch}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
*
*For logic simulation:
VA A 0 PULSE(3.3 0 0 1n 1n 1000n 2000n)
VB B 0 PULSE(3.3 0 0 1n 1n 500n 1000n)
*VC C 0 PULSE(3.3 0 0 1n 1n 250n 500n)
*VD D 0 PULSE(3.3 0 0 1n 1n 125n 250n)
*
.TRAN 0 2000n
.include Z:\MOS_model.txt
.END
